module name(
);
    logic a;
    wire b;

endmodule