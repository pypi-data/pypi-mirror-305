module ansi_module_d(
    input var logic a, b,
    output tri logic c,
    input wire d,
    inout e
);
    
endmodule