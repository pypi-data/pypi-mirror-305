module ansi_module_b;

  logic a;
  logic b;

endmodule
