module ansi_module_b (
  input var logic hej
);

  logic a;
  logic b;

endmodule
